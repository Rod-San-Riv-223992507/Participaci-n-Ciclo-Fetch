module MI(
    input [31:0] DirInst, 
    output reg [31:0] InstS
);

reg [31:0] MEM [0:31];  

initial begin
    
    MEM[0] = 32'b00000000000000000000000000000000;  
    MEM[1] = 32'b00000000000000000000000000000000;  
    MEM[2] = 32'b00000000000000000000000000000000;  
    MEM[3] = 32'b00000000000000000000000000000000;  
    MEM[4] = 32'b00000000000000000000000000000001;  
    MEM[5] = 32'b00000000000000000000000000000001;  
    MEM[6] = 32'b00000000000000000000000000000001;  
    MEM[7] = 32'b00000000000000000000000000000001;  
    MEM[8] = 32'b00000000000000000000000000000010;  
    MEM[9] = 32'b00000000000000000000000000000010;  
    MEM[10] = 32'b00000000000000000000000000000010;
    MEM[11] = 32'b00000000000000000000000000000010;
    MEM[12] = 32'b00000000000000000000000000000011;
    MEM[13] = 32'b00000000000000000000000000000011;
    MEM[14] = 32'b00000000000000000000000000000011;
    MEM[15] = 32'b00000000000000000000000000000011;
    
    
end

always @* begin
    InstS = MEM[DirInst];  
end

endmodule
